module MIPS(
    
)